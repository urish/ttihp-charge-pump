* NGSPICE file created from tt_um_urish_dickson_pump.ext - technology: ihp-sg13g2

.subckt tt_um_urish_dickson_pump VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2]
+ ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3]
+ uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3]
+ uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3]
+ uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3]
+ uo_out[4] uo_out[5] uo_out[6] uo_out[7] ua[0] ua[1] ua[2] ua[3]
X0 uo_out[7].t24 a_33768_28803.t6 nmos_diode_0/ntap1$1_0.well.t2 uo_out[7].t29 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X1 uo_out[7].t22 a_33768_28803.t6 nmos_diode_0/ntap1$1_0.well.t11 uo_out[7].t28 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X2 uo_out[7].t31 clk.t0 a_36767_28881# uo_out[7].t30 sg13_lv_nmos ad=0.1331p pd=1.12u as=0.1216p ps=1.02u w=0.64u l=0.13u
X3 nmos_diode_0/ntap1$1_0.well.t6 a_33768_28803.t6 VPWR.t7 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X4 sg13g2_and2_2_0.X.t2 nmos_diode_1/ntap1$1_0.well.t4 cap_cmim l=30u w=30u
X5 VPWR.t13 a_33768_28803.t6 nmos_diode_0/ntap1$1_0.well.t8 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X6 VPWR.t12 a_33768_28803.t6 nmos_diode_0/ntap1$1_0.well.t6 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X7 nmos_diode_3/ntap1$1_0.well.t2 nmos_diode_3/ntap1$1_0.well.t0 nmos_diode_2/ntap1$1_0.well.t0 nmos_diode_3/ntap1$1_0.well.t1 sg13_lv_nmos ad=4.08p pd=24.68u as=4.08p ps=24.68u w=12u l=0.13u
X8 VPWR.t11 a_33768_28803.t6 nmos_diode_0/ntap1$1_0.well.t4 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X9 uo_out[7].t27 a_33768_28803.t6 nmos_diode_0/ntap1$1_0.well.t0 uo_out[7].t26 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X10 a_33768_28803.t1 ena.t0 uo_out[7].t42 uo_out[7].t47 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X11 uo_out[7].t34 a_36673_28881# sg13g2_and2_2_0.X.t0 uo_out[7].t33 sg13_lv_nmos ad=0.2812p pd=2.24u as=0.1406p ps=1.12u w=0.74u l=0.13u
X12 VPWR.t14 a_33768_28803.t6 nmos_diode_0/ntap1$1_0.well.t14 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X13 a_33768_28803.t5 ena.t0 VPWR.t26 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X14 nmos_diode_2/ntap1$1_0.well.t3 nmos_diode_2/ntap1$1_0.well.t1 nmos_diode_1/ntap1$1_0.well.t0 nmos_diode_2/ntap1$1_0.well.t2 sg13_lv_nmos ad=4.08p pd=24.68u as=4.08p ps=24.68u w=12u l=0.13u
X15 nmos_diode_0/ntap1$1_0.well.t13 a_33768_28803.t6 uo_out[7].t6 uo_out[7].t25 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X16 nmos_diode_0/ntap1$1_0.well.t1 a_33768_28803.t6 uo_out[7].t24 uo_out[7].t23 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X17 nmos_diode_0/ntap1$1_0.well.t10 a_33768_28803.t6 uo_out[7].t22 uo_out[7].t21 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X18 nmos_diode_0/ntap1$1_0.well.t7 a_33768_28803.t6 VPWR.t13 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X19 nmos_diode_0/ntap1$1_0.well.t5 a_33768_28803.t6 VPWR.t12 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X20 sg13g2_inv_1_0.Y clk.t1 uo_out[7].t36 uo_out[7].t35 sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X21 nmos_diode_0/ntap1$1_0.well.t18 nmos_diode_0/ntap1$1_0.well.t16 nmos_diode_3/ntap1$1_0.well.t4 nmos_diode_0/ntap1$1_0.well.t17 sg13_lv_nmos ad=4.08p pd=24.68u as=4.08p ps=24.68u w=12u l=0.13u
X22 nmos_diode_0/ntap1$1_0.well.t3 a_33768_28803.t6 VPWR.t11 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X23 a_36097_28881# ena.t1 VPWR.t23 VPWR.t0 sg13_lv_pmos ad=0.1596p pd=1.22u as=0.2856p ps=2.36u w=0.84u l=0.13u
X24 nmos_diode_0/ntap1$1_0.well.t9 a_33768_28803.t6 uo_out[7].t20 uo_out[7].t19 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X25 uo_out[7].t44 ena.t0 a_33768_28803.t1 uo_out[7].t46 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X26 ua[0].t1 uo_out[7].t0 cap_cmim l=30u w=30u
X27 sg13g2_and2_2_0.X.t3 nmos_diode_3/ntap1$1_0.well.t3 cap_cmim l=30u w=30u
X28 uo_out[7].t12 a_33768_28803.t6 nmos_diode_0/ntap1$1_0.well.t9 uo_out[7].t18 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X29 uo_out[7].t10 a_33768_28803.t6 nmos_diode_0/ntap1$1_0.well.t13 uo_out[7].t17 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X30 a_33768_28803.t2 ena.t0 uo_out[7].t27 uo_out[7].t45 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X31 sg13g2_and2_2_1.X.t1 a_36097_28881# VPWR.t2 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.1918p ps=1.5u w=1.12u l=0.13u
X32 sg13g2_and2_2_1.X.t2 nmos_diode_2/ntap1$1_0.well.t4 cap_cmim l=30u w=30u
X33 nmos_diode_0/ntap1$1_0.well.t15 a_33768_28803.t6 VPWR.t10 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3976p ps=2.95u w=1.12u l=0.13u
X34 VPWR.t27 ena.t0 a_33768_28803.t5 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X35 a_36673_28881# ena.t2 VPWR.t24 VPWR.t0 sg13_lv_pmos ad=0.1596p pd=1.22u as=0.2856p ps=2.36u w=0.84u l=0.13u
X36 a_36191_28881# ena.t1 a_36097_28881# uo_out[7].t37 sg13_lv_nmos ad=0.1216p pd=1.02u as=0.2176p ps=1.96u w=0.64u l=0.13u
X37 VPWR.t4 a_33768_28803.t6 nmos_diode_0/ntap1$1_0.well.t15 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X38 VPWR.t3 a_33768_28803.t6 nmos_diode_0/ntap1$1_0.well.t5 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X39 VPWR.t1 a_36097_28881# sg13g2_and2_2_1.X.t1 VPWR.t0 sg13_lv_pmos ad=0.4256p pd=3u as=0.2128p ps=1.5u w=1.12u l=0.13u
X40 a_33768_28803.t3 ena.t0 VPWR.t14 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X41 uo_out[7].t14 a_33768_28803.t6 nmos_diode_0/ntap1$1_0.well.t1 uo_out[7].t16 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X42 uo_out[7].t8 a_33768_28803.t6 nmos_diode_0/ntap1$1_0.well.t10 uo_out[7].t15 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X43 sg13g2_and2_2_0.X.t1 a_36673_28881# VPWR.t19 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.1918p ps=1.5u w=1.12u l=0.13u
X44 sg13g2_inv_1_0.Y clk.t1 VPWR.t20 VPWR.t0 sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X45 nmos_diode_0/ntap1$1_0.well.t11 a_33768_28803.t6 uo_out[7].t14 uo_out[7].t13 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X46 a_36767_28881# ena.t2 a_36673_28881# uo_out[7].t38 sg13_lv_nmos ad=0.1216p pd=1.02u as=0.2176p ps=1.96u w=0.64u l=0.13u
X47 VPWR.t7 a_33768_28803.t6 nmos_diode_0/ntap1$1_0.well.t7 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X48 VPWR.t5 a_33768_28803.t6 nmos_diode_0/ntap1$1_0.well.t3 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X49 VPWR.t2 sg13g2_inv_1_0.Y a_36097_28881# VPWR.t0 sg13_lv_pmos ad=0.1918p pd=1.5u as=0.1596p ps=1.22u w=0.84u l=0.13u
X50 a_33768_28803.t0 ena.t0 uo_out[7].t44 uo_out[7].t43 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X51 nmos_diode_1/ntap1$1_0.well.t3 nmos_diode_1/ntap1$1_0.well.t1 ua[0].t0 nmos_diode_1/ntap1$1_0.well.t2 sg13_lv_nmos ad=4.08p pd=24.68u as=4.08p ps=24.68u w=12u l=0.13u
X52 nmos_diode_0/ntap1$1_0.well.t8 a_33768_28803.t6 VPWR.t5 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X53 sg13g2_and2_2_1.X.t0 a_36097_28881# uo_out[7].t4 uo_out[7].t3 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1331p ps=1.12u w=0.74u l=0.13u
X54 nmos_diode_0/ntap1$1_0.well.t2 a_33768_28803.t6 uo_out[7].t12 uo_out[7].t11 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X55 nmos_diode_0/ntap1$1_0.well.t0 a_33768_28803.t6 uo_out[7].t10 uo_out[7].t9 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X56 uo_out[7].t42 ena.t0 a_33768_28803.t2 uo_out[7].t41 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X57 uo_out[7].t40 ena.t0 a_33768_28803.t0 uo_out[7].t39 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
X58 uo_out[7].t2 a_36097_28881# sg13g2_and2_2_1.X.t0 uo_out[7].t1 sg13_lv_nmos ad=0.2812p pd=2.24u as=0.1406p ps=1.12u w=0.74u l=0.13u
X59 a_33768_28803.t4 ena.t0 VPWR.t27 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X60 VPWR.t19 clk.t0 a_36673_28881# VPWR.t0 sg13_lv_pmos ad=0.1918p pd=1.5u as=0.1596p ps=1.22u w=0.84u l=0.13u
X61 VPWR.t21 a_36673_28881# sg13g2_and2_2_0.X.t1 VPWR.t0 sg13_lv_pmos ad=0.4256p pd=3u as=0.2128p ps=1.5u w=1.12u l=0.13u
X62 uo_out[7].t4 sg13g2_inv_1_0.Y a_36191_28881# uo_out[7].t48 sg13_lv_nmos ad=0.1331p pd=1.12u as=0.1216p ps=1.02u w=0.64u l=0.13u
X63 nmos_diode_0/ntap1$1_0.well.t4 a_33768_28803.t6 VPWR.t4 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X64 nmos_diode_0/ntap1$1_0.well.t14 a_33768_28803.t6 VPWR.t3 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X65 VPWR.t26 ena.t0 a_33768_28803.t3 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X66 VPWR.t25 ena.t0 a_33768_28803.t4 VPWR.t0 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X67 nmos_diode_0/ntap1$1_0.well.t12 a_33768_28803.t6 uo_out[7].t8 uo_out[7].t7 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X68 sg13g2_and2_2_0.X.t0 a_36673_28881# uo_out[7].t31 uo_out[7].t32 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1331p ps=1.12u w=0.74u l=0.13u
X69 uo_out[7].t6 a_33768_28803.t6 nmos_diode_0/ntap1$1_0.well.t12 uo_out[7].t5 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
R0 a_33768_28803.n0 a_33768_28803.t6 13.4782
R1 a_33768_28803.n2 a_33768_28803.t0 9.07551
R2 a_33768_28803.n2 a_33768_28803.t1 8.58375
R3 a_33768_28803.n0 a_33768_28803.t2 8.58375
R4 a_33768_28803.n1 a_33768_28803.t4 6.26103
R5 a_33768_28803.n1 a_33768_28803.t3 5.7697
R6 a_33768_28803.t5 a_33768_28803.n1 5.76827
R7 a_33768_28803.n1 a_33768_28803.n0 1.0076
R8 a_33768_28803.n0 a_33768_28803.n2 0.929029
R9 nmos_diode_0/ntap1$1_0.well.n0 sg13g2_buf_16_0.X 18.7456
R10 nmos_diode_0/ntap1$1_0.well.n17 nmos_diode_0/ntap1$1_0.well.t16 15.0005
R11 nmos_diode_0/ntap1$1_0.well.n6 nmos_diode_0/ntap1$1_0.well.n4 9.43274
R12 nmos_diode_0/ntap1$1_0.well.n15 nmos_diode_0/ntap1$1_0.well.t2 9.0741
R13 nmos_diode_0/ntap1$1_0.well.n13 nmos_diode_0/ntap1$1_0.well.t1 9.0741
R14 nmos_diode_0/ntap1$1_0.well.n11 nmos_diode_0/ntap1$1_0.well.t11 9.0741
R15 nmos_diode_0/ntap1$1_0.well.n9 nmos_diode_0/ntap1$1_0.well.t10 9.0741
R16 nmos_diode_0/ntap1$1_0.well.n7 nmos_diode_0/ntap1$1_0.well.t12 9.0741
R17 nmos_diode_0/ntap1$1_0.well.n5 nmos_diode_0/ntap1$1_0.well.t13 9.0741
R18 nmos_diode_0/ntap1$1_0.well.n4 nmos_diode_0/ntap1$1_0.well.t0 9.0741
R19 nmos_diode_0/ntap1$1_0.well.n2 nmos_diode_0/ntap1$1_0.well.t9 9.0741
R20 nmos_diode_0/ntap1$1_0.well.n3 nmos_diode_0/ntap1$1_0.well.n2 9.04056
R21 nmos_diode_0/ntap1$1_0.well.n16 nmos_diode_0/ntap1$1_0.well.n15 9.04056
R22 nmos_diode_0/ntap1$1_0.well.n14 nmos_diode_0/ntap1$1_0.well.n13 9.04056
R23 nmos_diode_0/ntap1$1_0.well.n12 nmos_diode_0/ntap1$1_0.well.n11 9.04056
R24 nmos_diode_0/ntap1$1_0.well.n10 nmos_diode_0/ntap1$1_0.well.n9 9.04056
R25 nmos_diode_0/ntap1$1_0.well.n8 nmos_diode_0/ntap1$1_0.well.n7 9.04056
R26 nmos_diode_0/ntap1$1_0.well.n6 nmos_diode_0/ntap1$1_0.well.n5 9.04056
R27 nmos_diode_0/ntap1$1_0.well.n1 nmos_diode_0/ntap1$1_0.well.t17 5129.68
R28 nmos_diode_0/ntap1$1_0.well.n1 nmos_diode_0/ntap1$1_0.well.n0 0.0328461
R29 nmos_diode_0/ntap1$1_0.well.n2 nmos_diode_0/ntap1$1_0.well.t15 5.67875
R30 nmos_diode_0/ntap1$1_0.well.n15 nmos_diode_0/ntap1$1_0.well.t4 5.67831
R31 nmos_diode_0/ntap1$1_0.well.n13 nmos_diode_0/ntap1$1_0.well.t3 5.67831
R32 nmos_diode_0/ntap1$1_0.well.n11 nmos_diode_0/ntap1$1_0.well.t8 5.67831
R33 nmos_diode_0/ntap1$1_0.well.n9 nmos_diode_0/ntap1$1_0.well.t7 5.67831
R34 nmos_diode_0/ntap1$1_0.well.n7 nmos_diode_0/ntap1$1_0.well.t6 5.67831
R35 nmos_diode_0/ntap1$1_0.well.n5 nmos_diode_0/ntap1$1_0.well.t5 5.67831
R36 nmos_diode_0/ntap1$1_0.well.n4 nmos_diode_0/ntap1$1_0.well.t14 5.67831
R37 nmos_diode_0/ntap1$1_1.well nmos_diode_0/ntap1$1_0.well.n1 2.38457
R38 nmos_diode_0/ntap1$1_0.well.n17 nmos_diode_0/ntap1$1_0.well.t18 2.2081
R39 nmos_diode_0/ntap1$1_0.well.n10 nmos_diode_0/ntap1$1_0.well.n8 0.392674
R40 nmos_diode_0/ntap1$1_0.well.n12 nmos_diode_0/ntap1$1_0.well.n10 0.390761
R41 nmos_diode_0/ntap1$1_0.well.n14 nmos_diode_0/ntap1$1_0.well.n12 0.390761
R42 nmos_diode_0/ntap1$1_0.well.n16 nmos_diode_0/ntap1$1_0.well.n14 0.390761
R43 nmos_diode_0/ntap1$1_0.well.n8 nmos_diode_0/ntap1$1_0.well.n6 0.388848
R44 nmos_diode_0/ntap1$1_0.well.n0 nmos_diode_0/ntap1$1_0.well.n17 0.242882
R45 sg13g2_buf_16_0.X nmos_diode_0/ntap1$1_0.well.n3 0.143978
R46 nmos_diode_0/ntap1$1_0.well.n3 sg13g2_buf_16_0.X 0.0598043
R47 sg13g2_buf_16_0.X nmos_diode_0/ntap1$1_0.well.n16 0.0559783
R48 uo_out[7].t19 uo_out[7].n39 25.3211
R49 uo_out[7].n39 uo_out[7].t35 23.3603
R50 uo_out[7].n72 uo_out[7].t34 17.358
R51 uo_out[7].n71 uo_out[7].t31 17.358
R52 uo_out[7].n67 uo_out[7].t2 17.358
R53 uo_out[7].n66 uo_out[7].t4 17.358
R54 uo_out[7].n60 uo_out[7].t44 17.2861
R55 uo_out[7].n58 uo_out[7].t42 17.2861
R56 uo_out[7].n55 uo_out[7].t27 17.2807
R57 uo_out[7].n76 uo_out[7].n75 17.0005
R58 uo_out[7].n75 uo_out[7].n40 17.0005
R59 uo_out[7].n75 uo_out[7].n36 17.0005
R60 uo_out[7].n75 uo_out[7].n42 17.0005
R61 uo_out[7].n75 uo_out[7].n31 17.0005
R62 uo_out[7].n75 uo_out[7].n43 17.0005
R63 uo_out[7].n75 uo_out[7].n28 17.0005
R64 uo_out[7].n75 uo_out[7].n44 17.0005
R65 uo_out[7].n75 uo_out[7].n26 17.0005
R66 uo_out[7].n75 uo_out[7].n45 17.0005
R67 uo_out[7].n75 uo_out[7].n25 17.0005
R68 uo_out[7].n75 uo_out[7].n48 17.0005
R69 uo_out[7].n75 uo_out[7].n24 17.0005
R70 uo_out[7].n75 uo_out[7].n51 17.0005
R71 uo_out[7].n75 uo_out[7].n23 17.0005
R72 uo_out[7].n75 uo_out[7].n54 17.0005
R73 uo_out[7].n75 uo_out[7].n22 17.0005
R74 uo_out[7].n75 uo_out[7].n57 17.0005
R75 uo_out[7].n75 uo_out[7].n20 17.0005
R76 uo_out[7].n75 uo_out[7].n63 17.0005
R77 uo_out[7].n75 uo_out[7].n19 17.0005
R78 uo_out[7].n75 uo_out[7].n17 17.0005
R79 uo_out[7].n75 uo_out[7].n65 17.0005
R80 uo_out[7].n75 uo_out[7].n15 17.0005
R81 uo_out[7].n75 uo_out[7].n13 17.0005
R82 uo_out[7].n75 uo_out[7].n70 17.0005
R83 uo_out[7].n75 uo_out[7].n11 17.0005
R84 uo_out[7].t33 uo_out[7].n10 16.1677
R85 uo_out[7].t1 uo_out[7].n14 13.7435
R86 uo_out[7].t39 uo_out[7].n18 12.1956
R87 uo_out[7].n14 uo_out[7].t38 11.886
R88 uo_out[7].n18 uo_out[7].t37 11.886
R89 uo_out[7].t35 uo_out[7].n10 9.76892
R90 uo_out[7].t46 uo_out[7].n20 9.59769
R91 uo_out[7].n57 uo_out[7].t47 9.59769
R92 uo_out[7].n42 uo_out[7].t29 9.59769
R93 uo_out[7].t11 uo_out[7].n36 9.59769
R94 uo_out[7].n70 uo_out[7].t32 9.28811
R95 uo_out[7].n65 uo_out[7].t3 9.28811
R96 uo_out[7].n95 uo_out[7].n94 9.04683
R97 uo_out[7].n80 uo_out[7].n79 9.04679
R98 uo_out[7].n79 uo_out[7].n78 9.0005
R99 uo_out[7].n83 uo_out[7].n82 9.0005
R100 uo_out[7].n84 uo_out[7].n8 9.0005
R101 uo_out[7].n86 uo_out[7].n85 9.0005
R102 uo_out[7].n4 uo_out[7].n3 9.0005
R103 uo_out[7].n93 uo_out[7].n92 9.0005
R104 uo_out[7].n82 uo_out[7].n81 9.0005
R105 uo_out[7].n8 uo_out[7].n7 9.0005
R106 uo_out[7].n87 uo_out[7].n86 9.0005
R107 uo_out[7].n5 uo_out[7].n4 9.0005
R108 uo_out[7].n92 uo_out[7].n91 9.0005
R109 uo_out[7].n2 uo_out[7].n1 9.0005
R110 uo_out[7].n7 uo_out[7].n6 9.0005
R111 uo_out[7].n88 uo_out[7].n87 9.0005
R112 uo_out[7].n89 uo_out[7].n5 9.0005
R113 uo_out[7].n91 uo_out[7].n90 9.0005
R114 uo_out[7].n1 uo_out[7].n0 9.0005
R115 uo_out[7].n96 uo_out[7].n95 9.0005
R116 uo_out[7].n63 uo_out[7].t43 8.97852
R117 uo_out[7].t41 uo_out[7].n22 8.97852
R118 uo_out[7].t23 uo_out[7].n31 8.97852
R119 uo_out[7].n40 uo_out[7].t18 8.97852
R120 uo_out[7].n74 uo_out[7].t36 8.76703
R121 uo_out[7].n52 uo_out[7].t10 8.76678
R122 uo_out[7].n46 uo_out[7].t8 8.76678
R123 uo_out[7].n29 uo_out[7].t22 8.76678
R124 uo_out[7].n34 uo_out[7].t24 8.76678
R125 uo_out[7].n37 uo_out[7].t12 8.76678
R126 uo_out[7].n9 uo_out[7].t20 8.76678
R127 uo_out[7].n61 uo_out[7].t40 8.76312
R128 uo_out[7].n49 uo_out[7].t6 8.75736
R129 uo_out[7].n32 uo_out[7].t14 8.75736
R130 uo_out[7].t30 uo_out[7].n13 8.66893
R131 uo_out[7].t48 uo_out[7].n17 8.66893
R132 uo_out[7].n75 uo_out[7].n38 8.47111
R133 uo_out[7].n75 uo_out[7].n35 8.47111
R134 uo_out[7].n75 uo_out[7].n33 8.47111
R135 uo_out[7].n75 uo_out[7].n30 8.47111
R136 uo_out[7].n75 uo_out[7].n27 8.47111
R137 uo_out[7].n75 uo_out[7].n50 8.47111
R138 uo_out[7].n75 uo_out[7].n53 8.47111
R139 uo_out[7].n75 uo_out[7].n56 8.47111
R140 uo_out[7].n75 uo_out[7].n59 8.47111
R141 uo_out[7].n75 uo_out[7].n62 8.47111
R142 uo_out[7].n75 uo_out[7].n68 8.47111
R143 uo_out[7].n75 uo_out[7].n73 8.47111
R144 uo_out[7].n54 uo_out[7].t45 8.35935
R145 uo_out[7].n43 uo_out[7].t16 8.35935
R146 uo_out[7].t26 uo_out[7].n23 7.74017
R147 uo_out[7].t13 uo_out[7].n28 7.74017
R148 uo_out[7].n51 uo_out[7].t9 7.121
R149 uo_out[7].n44 uo_out[7].t28 7.121
R150 uo_out[7].n75 uo_out[7].n41 6.58313
R151 uo_out[7].n75 uo_out[7].n21 6.58313
R152 uo_out[7].n75 uo_out[7].n18 6.58313
R153 uo_out[7].n75 uo_out[7].n16 6.58313
R154 uo_out[7].n75 uo_out[7].n14 6.58313
R155 uo_out[7].n75 uo_out[7].n12 6.58313
R156 uo_out[7].t17 uo_out[7].n24 6.50182
R157 uo_out[7].t21 uo_out[7].n26 6.50182
R158 uo_out[7].n97 uo_out[7].n96 6.28223
R159 uo_out[7].n48 uo_out[7].t25 5.88265
R160 uo_out[7].n45 uo_out[7].t15 5.88265
R161 uo_out[7].n75 uo_out[7].n74 5.66845
R162 uo_out[7].n75 uo_out[7].n47 5.61485
R163 uo_out[7].n75 uo_out[7].n64 5.61485
R164 uo_out[7].n75 uo_out[7].n69 5.61485
R165 uo_out[7].t5 uo_out[7].n25 5.26348
R166 uo_out[7].t7 uo_out[7].n25 5.26348
R167 uo_out[7].n48 uo_out[7].t5 4.6443
R168 uo_out[7].n45 uo_out[7].t7 4.6443
R169 uo_out[7].n94 uo_out[7].n93 4.59267
R170 uo_out[7].n80 uo_out[7].n6 4.56979
R171 uo_out[7].t32 uo_out[7].n12 4.45592
R172 uo_out[7].t3 uo_out[7].n16 4.45592
R173 uio_oe[7] uo_out[7].n116 4.2409
R174 uo_out[7].n21 uo_out[7].t46 4.14633
R175 uo_out[7].t47 uo_out[7].n21 4.14633
R176 uo_out[7].t29 uo_out[7].n41 4.14633
R177 uo_out[7].n41 uo_out[7].t11 4.14633
R178 uo_out[7].t25 uo_out[7].n24 4.02513
R179 uo_out[7].t15 uo_out[7].n26 4.02513
R180 uo_out[7].n16 uo_out[7].t1 3.83675
R181 uo_out[7].n12 uo_out[7].t33 3.83675
R182 uo_out[7].n51 uo_out[7].t17 3.40596
R183 uo_out[7].n44 uo_out[7].t21 3.40596
R184 uo_out[7].n116 VGND 3.2345
R185 uo_out[7].n114 VGND 3.1465
R186 uo_out[7].n75 uo_out[7].n10 2.99906
R187 uo_out[7].t9 uo_out[7].n23 2.78678
R188 uo_out[7].t28 uo_out[7].n28 2.78678
R189 uo_out[7].n78 uo_out[7].n77 2.50974
R190 uo_out[7].n54 uo_out[7].t26 2.16761
R191 uo_out[7].n43 uo_out[7].t13 2.16761
R192 uo_out[7].t38 uo_out[7].n13 1.85802
R193 uo_out[7].t37 uo_out[7].n17 1.85802
R194 uo_out[7].n63 uo_out[7].t39 1.54843
R195 uo_out[7].t45 uo_out[7].n22 1.54843
R196 uo_out[7].t16 uo_out[7].n31 1.54843
R197 uo_out[7].n40 uo_out[7].t19 1.54843
R198 uo_out[7].n70 uo_out[7].t30 1.23885
R199 uo_out[7].n65 uo_out[7].t48 1.23885
R200 uo_out[7].t43 uo_out[7].n20 0.929261
R201 uo_out[7].n57 uo_out[7].t41 0.929261
R202 uo_out[7].n42 uo_out[7].t23 0.929261
R203 uo_out[7].t18 uo_out[7].n36 0.929261
R204 uo_out[7].n114 VGND 0.851816
R205 uo_out[7].n99 uo_out[1] 0.5417
R206 uo_out[7].n100 uo_out[2] 0.5417
R207 uo_out[7].n101 uo_out[3] 0.5417
R208 uo_out[7].n102 uo_out[4] 0.5417
R209 uo_out[7].n103 uo_out[5] 0.5417
R210 uo_out[7].n104 uo_out[6] 0.5417
R211 uo_out[7].n105 uo_out[7] 0.5417
R212 uo_out[7].n106 uio_out[0] 0.5417
R213 uo_out[7].n107 uio_out[1] 0.5417
R214 uo_out[7].n108 uio_out[2] 0.5417
R215 uo_out[7].n109 uio_out[3] 0.5417
R216 uo_out[7].n110 uio_out[4] 0.5417
R217 uo_out[7].n111 uio_out[5] 0.5417
R218 uo_out[7].n112 uio_out[6] 0.5417
R219 uo_out[7].n113 uio_out[7] 0.5417
R220 uio_oe[0] uo_out[7].n123 0.5417
R221 uio_oe[1] uo_out[7].n122 0.5417
R222 uio_oe[2] uo_out[7].n121 0.5417
R223 uio_oe[3] uo_out[7].n120 0.5417
R224 uio_oe[4] uo_out[7].n119 0.5417
R225 uio_oe[5] uo_out[7].n118 0.5417
R226 uio_oe[6] uo_out[7].n117 0.5417
R227 uo_out[7].n98 uo_out[7].n97 0.540233
R228 uo_out[7].n69 uo_out[7] 0.180825
R229 uo_out[7].n64 uo_out[7] 0.180825
R230 uo_out[7].n50 uo_out[7].n49 0.173289
R231 uo_out[7].n46 uo_out[7].n27 0.173289
R232 uo_out[7].n71 uo_out[7].n69 0.169236
R233 uo_out[7].n66 uo_out[7].n64 0.169236
R234 uo_out[7].n53 uo_out[7].n52 0.158289
R235 uo_out[7].n30 uo_out[7].n29 0.158289
R236 uo_out[7].n62 uo_out[7].n61 0.143289
R237 uo_out[7].n56 uo_out[7].n55 0.143289
R238 uo_out[7].n33 uo_out[7].n32 0.143289
R239 uo_out[7].n38 uo_out[7].n9 0.143289
R240 uo_out[7].n73 uo_out[7].n71 0.132039
R241 uo_out[7].n68 uo_out[7].n66 0.132039
R242 uo_out[7].n47 uo_out[7].n46 0.128325
R243 uo_out[7].n60 uo_out[7].n59 0.128289
R244 uo_out[7].n59 uo_out[7].n58 0.128289
R245 uo_out[7].n35 uo_out[7].n34 0.128289
R246 uo_out[7].n37 uo_out[7].n35 0.128289
R247 uo_out[7].n49 uo_out[7].n47 0.127986
R248 uo_out[7].n74 uo_out[7] 0.126449
R249 uo_out[7].n73 uo_out[7].n72 0.124539
R250 uo_out[7].n68 uo_out[7].n67 0.124539
R251 uo_out[7].n62 uo_out[7].n60 0.113289
R252 uo_out[7].n58 uo_out[7].n56 0.113289
R253 uo_out[7].n34 uo_out[7].n33 0.113289
R254 uo_out[7].n38 uo_out[7].n37 0.113289
R255 uo_out[7].n55 uo_out[7].n53 0.098289
R256 uo_out[7].n32 uo_out[7].n30 0.098289
R257 uo_out[7].n83 uo_out[7].n78 0.0921667
R258 uo_out[7].n84 uo_out[7].n83 0.0921667
R259 uo_out[7].n85 uo_out[7].n84 0.0921667
R260 uo_out[7].n85 uo_out[7].n3 0.0921667
R261 uo_out[7].n93 uo_out[7].n3 0.0921667
R262 uo_out[7].n82 uo_out[7].n79 0.0921667
R263 uo_out[7].n82 uo_out[7].n8 0.0921667
R264 uo_out[7].n86 uo_out[7].n8 0.0921667
R265 uo_out[7].n86 uo_out[7].n4 0.0921667
R266 uo_out[7].n92 uo_out[7].n4 0.0921667
R267 uo_out[7].n92 uo_out[7].n2 0.0921667
R268 uo_out[7].n81 uo_out[7].n7 0.0921667
R269 uo_out[7].n87 uo_out[7].n7 0.0921667
R270 uo_out[7].n87 uo_out[7].n5 0.0921667
R271 uo_out[7].n91 uo_out[7].n5 0.0921667
R272 uo_out[7].n91 uo_out[7].n1 0.0921667
R273 uo_out[7].n95 uo_out[7].n1 0.0921667
R274 uo_out[7].n52 uo_out[7].n50 0.083289
R275 uo_out[7].n29 uo_out[7].n27 0.083289
R276 uo_out[7].n88 uo_out[7].n6 0.0738333
R277 uo_out[7].n89 uo_out[7].n88 0.0738333
R278 uo_out[7].n90 uo_out[7].n89 0.0738333
R279 uo_out[7].n90 uo_out[7].n0 0.0738333
R280 uo_out[7].n96 uo_out[7].n0 0.0738333
R281 uo_out[7] uo_out[7].n11 0.0605
R282 uo_out[7] uo_out[7].n15 0.0605
R283 uo_out[7] uo_out[7].n19 0.0605
R284 uo_out[7].n77 uo_out[7].n76 0.0591035
R285 uo_out[7].n72 uo_out[7].n11 0.05675
R286 uo_out[7].n67 uo_out[7].n15 0.05675
R287 uo_out[7].n81 uo_out[7].n80 0.046417
R288 uo_out[7].n94 uo_out[7].n2 0.0463712
R289 uo_out[7].n115 uo_out[7].t0 0.0445
R290 uo_out[7].n61 uo_out[7].n19 0.038
R291 uo_out[7].n76 uo_out[7].n9 0.038
R292 uo_out[1] uo_out[7].n98 0.0225
R293 uo_out[2] uo_out[7].n99 0.0225
R294 uo_out[3] uo_out[7].n100 0.0225
R295 uo_out[4] uo_out[7].n101 0.0225
R296 uo_out[5] uo_out[7].n102 0.0225
R297 uo_out[6] uo_out[7].n103 0.0225
R298 uo_out[7] uo_out[7].n104 0.0225
R299 uio_out[0] uo_out[7].n105 0.0225
R300 uio_out[1] uo_out[7].n106 0.0225
R301 uio_out[2] uo_out[7].n107 0.0225
R302 uio_out[3] uo_out[7].n108 0.0225
R303 uio_out[4] uo_out[7].n109 0.0225
R304 uio_out[5] uo_out[7].n110 0.0225
R305 uio_out[6] uo_out[7].n111 0.0225
R306 uio_out[7] uo_out[7].n112 0.0225
R307 uio_oe[0] uo_out[7].n113 0.0225
R308 uo_out[7].n123 uio_oe[1] 0.0225
R309 uo_out[7].n122 uio_oe[2] 0.0225
R310 uo_out[7].n121 uio_oe[3] 0.0225
R311 uo_out[7].n120 uio_oe[4] 0.0225
R312 uo_out[7].n119 uio_oe[5] 0.0225
R313 uo_out[7].n118 uio_oe[6] 0.0225
R314 uo_out[7].n117 uio_oe[7] 0.0225
R315 uo_out[7].n75 uo_out[7].n39 0.0203952
R316 uo_out[7].n98 uo_out[1] 0.0155
R317 uo_out[7].n99 uo_out[2] 0.0155
R318 uo_out[7].n100 uo_out[3] 0.0155
R319 uo_out[7].n101 uo_out[4] 0.0155
R320 uo_out[7].n102 uo_out[5] 0.0155
R321 uo_out[7].n103 uo_out[6] 0.0155
R322 uo_out[7].n104 uo_out[7] 0.0155
R323 uo_out[7].n105 uio_out[0] 0.0155
R324 uo_out[7].n106 uio_out[1] 0.0155
R325 uo_out[7].n107 uio_out[2] 0.0155
R326 uo_out[7].n108 uio_out[3] 0.0155
R327 uo_out[7].n109 uio_out[4] 0.0155
R328 uo_out[7].n110 uio_out[5] 0.0155
R329 uo_out[7].n111 uio_out[6] 0.0155
R330 uo_out[7].n112 uio_out[7] 0.0155
R331 uo_out[7].n113 uio_oe[0] 0.0155
R332 uo_out[7].n123 uio_oe[1] 0.0155
R333 uo_out[7].n122 uio_oe[2] 0.0155
R334 uo_out[7].n121 uio_oe[3] 0.0155
R335 uo_out[7].n120 uio_oe[4] 0.0155
R336 uo_out[7].n119 uio_oe[5] 0.0155
R337 uo_out[7].n118 uio_oe[6] 0.0155
R338 uo_out[7].n117 uio_oe[7] 0.0155
R339 uo_out[7].n116 uo_out[7].n115 0.0124065
R340 uo_out[7].n115 uo_out[7].n114 0.0124065
R341 uo_out[7].n77 uo_out[7] 0.00285354
R342 uo_out[7].n97 uo_out[0] 0.00196667
R343 clk.n1 clk 29.7446
R344 clk.n0 clk.t0 15.0287
R345 clk.n1 clk.n0 9.6781
R346 clk.n2 clk.n1 9.01476
R347 clk.n2 clk.t1 7.50757
R348 clk clk.n2 0.0571086
R349 clk.n0 clk 0.0569103
R350 VPWR.n155 VPWR.n154 17.0005
R351 VPWR.n154 VPWR.n14 17.0005
R352 VPWR.n154 VPWR.n19 17.0005
R353 VPWR.n154 VPWR.n13 17.0005
R354 VPWR.n154 VPWR.n25 17.0005
R355 VPWR.n154 VPWR.n153 17.0005
R356 VPWR.n113 VPWR.n67 9.05107
R357 VPWR.n150 VPWR.n149 9.051
R358 VPWR.n117 VPWR.n67 9.05072
R359 VPWR.n112 VPWR.n69 9.0005
R360 VPWR.n111 VPWR.n110 9.0005
R361 VPWR.n109 VPWR.n70 9.0005
R362 VPWR.n108 VPWR.n107 9.0005
R363 VPWR.n106 VPWR.n72 9.0005
R364 VPWR.n105 VPWR.n104 9.0005
R365 VPWR.n103 VPWR.n73 9.0005
R366 VPWR.n102 VPWR.n101 9.0005
R367 VPWR.n100 VPWR.n75 9.0005
R368 VPWR.n99 VPWR.n98 9.0005
R369 VPWR.n97 VPWR.n76 9.0005
R370 VPWR.n96 VPWR.n95 9.0005
R371 VPWR.n94 VPWR.n78 9.0005
R372 VPWR.n93 VPWR.n92 9.0005
R373 VPWR.n91 VPWR.n79 9.0005
R374 VPWR.n90 VPWR.n89 9.0005
R375 VPWR.n88 VPWR.n81 9.0005
R376 VPWR.n87 VPWR.n86 9.0005
R377 VPWR.n85 VPWR.n82 9.0005
R378 VPWR.n84 VPWR.n83 9.0005
R379 VPWR.n39 VPWR.n38 9.0005
R380 VPWR.n152 VPWR.n151 9.0005
R381 VPWR.n40 VPWR.n39 9.0005
R382 VPWR.n84 VPWR.n43 9.0005
R383 VPWR.n85 VPWR.n44 9.0005
R384 VPWR.n86 VPWR.n45 9.0005
R385 VPWR.n81 VPWR.n80 9.0005
R386 VPWR.n90 VPWR.n48 9.0005
R387 VPWR.n91 VPWR.n49 9.0005
R388 VPWR.n92 VPWR.n50 9.0005
R389 VPWR.n78 VPWR.n77 9.0005
R390 VPWR.n96 VPWR.n53 9.0005
R391 VPWR.n97 VPWR.n54 9.0005
R392 VPWR.n98 VPWR.n55 9.0005
R393 VPWR.n75 VPWR.n74 9.0005
R394 VPWR.n102 VPWR.n58 9.0005
R395 VPWR.n103 VPWR.n59 9.0005
R396 VPWR.n104 VPWR.n60 9.0005
R397 VPWR.n72 VPWR.n71 9.0005
R398 VPWR.n108 VPWR.n63 9.0005
R399 VPWR.n109 VPWR.n64 9.0005
R400 VPWR.n110 VPWR.n65 9.0005
R401 VPWR.n69 VPWR.n68 9.0005
R402 VPWR.n115 VPWR.n114 9.0005
R403 VPWR.n151 VPWR.n150 9.0005
R404 VPWR.n41 VPWR.n40 9.0005
R405 VPWR.n147 VPWR.n43 9.0005
R406 VPWR.n146 VPWR.n44 9.0005
R407 VPWR.n145 VPWR.n45 9.0005
R408 VPWR.n80 VPWR.n46 9.0005
R409 VPWR.n141 VPWR.n48 9.0005
R410 VPWR.n140 VPWR.n49 9.0005
R411 VPWR.n139 VPWR.n50 9.0005
R412 VPWR.n77 VPWR.n51 9.0005
R413 VPWR.n135 VPWR.n53 9.0005
R414 VPWR.n134 VPWR.n54 9.0005
R415 VPWR.n133 VPWR.n55 9.0005
R416 VPWR.n74 VPWR.n56 9.0005
R417 VPWR.n129 VPWR.n58 9.0005
R418 VPWR.n128 VPWR.n59 9.0005
R419 VPWR.n127 VPWR.n60 9.0005
R420 VPWR.n71 VPWR.n61 9.0005
R421 VPWR.n123 VPWR.n63 9.0005
R422 VPWR.n122 VPWR.n64 9.0005
R423 VPWR.n121 VPWR.n65 9.0005
R424 VPWR.n68 VPWR.n66 9.0005
R425 VPWR.n116 VPWR.n115 9.0005
R426 VPWR.n148 VPWR.n147 9.0005
R427 VPWR.n146 VPWR.n42 9.0005
R428 VPWR.n145 VPWR.n144 9.0005
R429 VPWR.n143 VPWR.n46 9.0005
R430 VPWR.n142 VPWR.n141 9.0005
R431 VPWR.n140 VPWR.n47 9.0005
R432 VPWR.n139 VPWR.n138 9.0005
R433 VPWR.n137 VPWR.n51 9.0005
R434 VPWR.n136 VPWR.n135 9.0005
R435 VPWR.n134 VPWR.n52 9.0005
R436 VPWR.n133 VPWR.n132 9.0005
R437 VPWR.n131 VPWR.n56 9.0005
R438 VPWR.n130 VPWR.n129 9.0005
R439 VPWR.n128 VPWR.n57 9.0005
R440 VPWR.n127 VPWR.n126 9.0005
R441 VPWR.n125 VPWR.n61 9.0005
R442 VPWR.n124 VPWR.n123 9.0005
R443 VPWR.n122 VPWR.n62 9.0005
R444 VPWR.n23 VPWR.t23 8.78204
R445 VPWR.n17 VPWR.t24 8.78204
R446 VPWR.n22 VPWR.t2 8.77677
R447 VPWR.n20 VPWR.t1 8.77677
R448 VPWR.n16 VPWR.t19 8.77677
R449 VPWR.n1 VPWR.t21 8.77677
R450 VPWR.n32 VPWR.t14 8.77315
R451 VPWR.n30 VPWR.t26 8.77315
R452 VPWR.n28 VPWR.t27 8.77315
R453 VPWR.n154 VPWR.n15 8.47111
R454 VPWR.n154 VPWR.n18 8.47111
R455 VPWR.n154 VPWR.n21 8.47111
R456 VPWR.n154 VPWR.n24 8.47111
R457 VPWR.n154 VPWR.n27 8.47111
R458 VPWR.n154 VPWR.n29 8.47111
R459 VPWR.n154 VPWR.n31 8.47111
R460 VPWR.n154 VPWR.n33 8.47111
R461 VPWR.n154 VPWR.n36 8.47111
R462 VPWR.n154 VPWR.n10 8.47111
R463 VPWR.n154 VPWR.n8 8.47111
R464 VPWR.n154 VPWR.n6 8.47111
R465 VPWR.n154 VPWR.n4 8.47111
R466 VPWR.n154 VPWR.n2 8.47111
R467 VPWR.n0 VPWR.t20 5.99762
R468 VPWR.n37 VPWR.t10 5.99168
R469 VPWR.n26 VPWR.t25 5.98924
R470 VPWR.n3 VPWR.t4 5.98777
R471 VPWR.n5 VPWR.t11 5.98777
R472 VPWR.n9 VPWR.t13 5.98777
R473 VPWR.n35 VPWR.t12 5.98777
R474 VPWR.n11 VPWR.t7 5.98658
R475 VPWR.n34 VPWR.t3 5.98658
R476 VPWR.n7 VPWR.t5 5.98588
R477 VPWR.n118 VPWR 5.7963
R478 VPWR.n154 VPWR.n0 5.66762
R479 VPWR.n154 VPWR.n12 5.61485
R480 VPWR.n113 VPWR.n112 4.63217
R481 VPWR.n149 VPWR.n148 4.601
R482 VPWR.n120 VPWR.n119 4.47614
R483 VPWR.n119 VPWR.n117 4.47614
R484 VPWR.n154 VPWR.t0 0.4255
R485 VPWR.n36 VPWR.n35 0.173289
R486 VPWR.n11 VPWR.n10 0.173289
R487 VPWR.n34 VPWR.n33 0.158289
R488 VPWR.n9 VPWR.n8 0.158289
R489 VPWR.n18 VPWR.n17 0.147039
R490 VPWR.n24 VPWR.n23 0.147039
R491 VPWR.n27 VPWR.n26 0.143289
R492 VPWR.n32 VPWR.n31 0.143289
R493 VPWR.n7 VPWR.n6 0.143289
R494 VPWR.n37 VPWR.n2 0.143289
R495 VPWR.n16 VPWR.n15 0.132039
R496 VPWR.n22 VPWR.n21 0.132039
R497 VPWR.n35 VPWR.n12 0.128325
R498 VPWR.n29 VPWR.n28 0.128289
R499 VPWR.n30 VPWR.n29 0.128289
R500 VPWR.n5 VPWR.n4 0.128289
R501 VPWR.n4 VPWR.n3 0.128289
R502 VPWR.n12 VPWR.n11 0.127986
R503 VPWR VPWR.n0 0.127277
R504 VPWR.n152 VPWR.n38 0.1255
R505 VPWR.n83 VPWR.n38 0.1255
R506 VPWR.n83 VPWR.n82 0.1255
R507 VPWR.n87 VPWR.n82 0.1255
R508 VPWR.n88 VPWR.n87 0.1255
R509 VPWR.n89 VPWR.n88 0.1255
R510 VPWR.n89 VPWR.n79 0.1255
R511 VPWR.n93 VPWR.n79 0.1255
R512 VPWR.n94 VPWR.n93 0.1255
R513 VPWR.n95 VPWR.n94 0.1255
R514 VPWR.n95 VPWR.n76 0.1255
R515 VPWR.n99 VPWR.n76 0.1255
R516 VPWR.n100 VPWR.n99 0.1255
R517 VPWR.n101 VPWR.n100 0.1255
R518 VPWR.n101 VPWR.n73 0.1255
R519 VPWR.n105 VPWR.n73 0.1255
R520 VPWR.n106 VPWR.n105 0.1255
R521 VPWR.n107 VPWR.n106 0.1255
R522 VPWR.n107 VPWR.n70 0.1255
R523 VPWR.n111 VPWR.n70 0.1255
R524 VPWR.n112 VPWR.n111 0.1255
R525 VPWR.n15 VPWR.n1 0.124539
R526 VPWR.n21 VPWR.n20 0.124539
R527 VPWR.n28 VPWR.n27 0.113289
R528 VPWR.n31 VPWR.n30 0.113289
R529 VPWR.n6 VPWR.n5 0.113289
R530 VPWR.n3 VPWR.n2 0.113289
R531 VPWR.n18 VPWR.n16 0.109539
R532 VPWR.n24 VPWR.n22 0.109539
R533 VPWR.n151 VPWR.n39 0.1005
R534 VPWR.n84 VPWR.n39 0.1005
R535 VPWR.n85 VPWR.n84 0.1005
R536 VPWR.n86 VPWR.n85 0.1005
R537 VPWR.n86 VPWR.n81 0.1005
R538 VPWR.n90 VPWR.n81 0.1005
R539 VPWR.n91 VPWR.n90 0.1005
R540 VPWR.n92 VPWR.n91 0.1005
R541 VPWR.n92 VPWR.n78 0.1005
R542 VPWR.n96 VPWR.n78 0.1005
R543 VPWR.n97 VPWR.n96 0.1005
R544 VPWR.n98 VPWR.n97 0.1005
R545 VPWR.n98 VPWR.n75 0.1005
R546 VPWR.n102 VPWR.n75 0.1005
R547 VPWR.n103 VPWR.n102 0.1005
R548 VPWR.n104 VPWR.n103 0.1005
R549 VPWR.n104 VPWR.n72 0.1005
R550 VPWR.n108 VPWR.n72 0.1005
R551 VPWR.n109 VPWR.n108 0.1005
R552 VPWR.n110 VPWR.n109 0.1005
R553 VPWR.n110 VPWR.n69 0.1005
R554 VPWR.n114 VPWR.n69 0.1005
R555 VPWR.n150 VPWR.n40 0.1005
R556 VPWR.n43 VPWR.n40 0.1005
R557 VPWR.n44 VPWR.n43 0.1005
R558 VPWR.n45 VPWR.n44 0.1005
R559 VPWR.n80 VPWR.n45 0.1005
R560 VPWR.n80 VPWR.n48 0.1005
R561 VPWR.n49 VPWR.n48 0.1005
R562 VPWR.n50 VPWR.n49 0.1005
R563 VPWR.n77 VPWR.n50 0.1005
R564 VPWR.n77 VPWR.n53 0.1005
R565 VPWR.n54 VPWR.n53 0.1005
R566 VPWR.n55 VPWR.n54 0.1005
R567 VPWR.n74 VPWR.n55 0.1005
R568 VPWR.n74 VPWR.n58 0.1005
R569 VPWR.n59 VPWR.n58 0.1005
R570 VPWR.n60 VPWR.n59 0.1005
R571 VPWR.n71 VPWR.n60 0.1005
R572 VPWR.n71 VPWR.n63 0.1005
R573 VPWR.n64 VPWR.n63 0.1005
R574 VPWR.n65 VPWR.n64 0.1005
R575 VPWR.n68 VPWR.n65 0.1005
R576 VPWR.n115 VPWR.n68 0.1005
R577 VPWR.n115 VPWR.n67 0.1005
R578 VPWR.n147 VPWR.n41 0.1005
R579 VPWR.n147 VPWR.n146 0.1005
R580 VPWR.n146 VPWR.n145 0.1005
R581 VPWR.n145 VPWR.n46 0.1005
R582 VPWR.n141 VPWR.n46 0.1005
R583 VPWR.n141 VPWR.n140 0.1005
R584 VPWR.n140 VPWR.n139 0.1005
R585 VPWR.n139 VPWR.n51 0.1005
R586 VPWR.n135 VPWR.n51 0.1005
R587 VPWR.n135 VPWR.n134 0.1005
R588 VPWR.n134 VPWR.n133 0.1005
R589 VPWR.n133 VPWR.n56 0.1005
R590 VPWR.n129 VPWR.n56 0.1005
R591 VPWR.n129 VPWR.n128 0.1005
R592 VPWR.n128 VPWR.n127 0.1005
R593 VPWR.n127 VPWR.n61 0.1005
R594 VPWR.n123 VPWR.n61 0.1005
R595 VPWR.n123 VPWR.n122 0.1005
R596 VPWR.n122 VPWR.n121 0.1005
R597 VPWR.n116 VPWR.n66 0.1005
R598 VPWR.n148 VPWR.n42 0.1005
R599 VPWR.n144 VPWR.n42 0.1005
R600 VPWR.n144 VPWR.n143 0.1005
R601 VPWR.n143 VPWR.n142 0.1005
R602 VPWR.n142 VPWR.n47 0.1005
R603 VPWR.n138 VPWR.n47 0.1005
R604 VPWR.n138 VPWR.n137 0.1005
R605 VPWR.n137 VPWR.n136 0.1005
R606 VPWR.n136 VPWR.n52 0.1005
R607 VPWR.n132 VPWR.n52 0.1005
R608 VPWR.n132 VPWR.n131 0.1005
R609 VPWR.n131 VPWR.n130 0.1005
R610 VPWR.n130 VPWR.n57 0.1005
R611 VPWR.n126 VPWR.n57 0.1005
R612 VPWR.n126 VPWR.n125 0.1005
R613 VPWR.n125 VPWR.n124 0.1005
R614 VPWR.n124 VPWR.n62 0.1005
R615 VPWR.n33 VPWR.n32 0.098289
R616 VPWR.n8 VPWR.n7 0.098289
R617 VPWR.n36 VPWR.n34 0.083289
R618 VPWR.n10 VPWR.n9 0.083289
R619 VPWR.n118 VPWR.n62 0.0685
R620 VPWR VPWR.n155 0.0605
R621 VPWR VPWR.n14 0.0605
R622 VPWR.n19 VPWR 0.0605
R623 VPWR VPWR.n13 0.0605
R624 VPWR.n25 VPWR 0.0605
R625 VPWR.n153 VPWR 0.0605
R626 VPWR.n155 VPWR.n1 0.05675
R627 VPWR.n20 VPWR.n19 0.05675
R628 VPWR VPWR.n152 0.0555
R629 VPWR.n121 VPWR.n120 0.0507238
R630 VPWR.n117 VPWR.n116 0.0507238
R631 VPWR.n120 VPWR.n66 0.0507238
R632 VPWR.n149 VPWR.n41 0.0504506
R633 VPWR.n114 VPWR.n113 0.0503827
R634 VPWR.n26 VPWR.n25 0.038
R635 VPWR.n153 VPWR.n37 0.038
R636 VPWR.n17 VPWR.n14 0.03425
R637 VPWR.n23 VPWR.n13 0.03425
R638 VPWR.n119 VPWR.n118 0.0007
R639 sg13g2_and2_2_0.X.n0 sg13g2_and2_2_0.X.t2 50.6368
R640 sg13g2_and2_2_0.X.n0 sg13g2_and2_2_0.X.t3 31.8635
R641 sg13g2_and2_2_0.X sg13g2_and2_2_0.X.n0 20.4337
R642 sg13g2_and2_2_0.X sg13g2_and2_2_0.X.t0 9.02933
R643 sg13g2_and2_2_0.X sg13g2_and2_2_0.X.t1 5.7736
R644 nmos_diode_1/ntap1$1_0.well.n2 nmos_diode_1/ntap1$1_0.well.t4 29.5591
R645 nmos_diode_1/ntap1$1_0.well.n3 nmos_diode_1/ntap1$1_0.well.t1 15.0005
R646 nmos_diode_1/ntap1$1_0.well.n0 nmos_diode_1/ntap1$1_0.well.n1 0.0328461
R647 nmos_diode_1/ntap1$1_0.well.t2 nmos_diode_1/ntap1$1_0.well.n1 5129.68
R648 nmos_diode_1/ntap1$1_0.well.n0 nmos_diode_1/ntap1$1_0.well.n2 7.10139
R649 nmos_diode_1/ntap1$1_0.well.n2 nmos_diode_1/ntap1$1_0.well.t0 6.54661
R650 nmos_diode_1/ntap1$1_0.well.n3 nmos_diode_1/ntap1$1_0.well.t3 2.2081
R651 nmos_diode_1/ntap1$1_1.well nmos_diode_1/ntap1$1_0.well.n0 2.35302
R652 nmos_diode_1/ntap1$1_0.well.n3 nmos_diode_1/ntap1$1_0.well.n1 0.275228
R653 nmos_diode_3/ntap1$1_0.well.n2 nmos_diode_3/ntap1$1_0.well.t3 29.7901
R654 nmos_diode_3/ntap1$1_0.well.n3 nmos_diode_3/ntap1$1_0.well.t0 15.0005
R655 nmos_diode_3/ntap1$1_0.well.n0 nmos_diode_3/ntap1$1_0.well.n1 0.0328461
R656 nmos_diode_3/ntap1$1_0.well.t1 nmos_diode_3/ntap1$1_0.well.n1 5129.68
R657 nmos_diode_3/ntap1$1_0.well.n0 nmos_diode_3/ntap1$1_0.well.n2 6.64037
R658 nmos_diode_3/ntap1$1_0.well.n2 nmos_diode_3/ntap1$1_0.well.t4 5.77135
R659 nmos_diode_3/ntap1$1_1.well nmos_diode_3/ntap1$1_0.well.n0 2.35223
R660 nmos_diode_3/ntap1$1_0.well.n3 nmos_diode_3/ntap1$1_0.well.t2 2.2081
R661 nmos_diode_3/ntap1$1_0.well.n3 nmos_diode_3/ntap1$1_0.well.n1 0.275228
R662 nmos_diode_2/ntap1$1_0.well.n2 nmos_diode_2/ntap1$1_0.well.t4 29.595
R663 nmos_diode_2/ntap1$1_0.well.n3 nmos_diode_2/ntap1$1_0.well.t1 15.0005
R664 nmos_diode_2/ntap1$1_0.well.n0 nmos_diode_2/ntap1$1_0.well.n1 0.0328461
R665 nmos_diode_2/ntap1$1_0.well.t2 nmos_diode_2/ntap1$1_0.well.n1 5129.68
R666 nmos_diode_2/ntap1$1_0.well.n0 nmos_diode_2/ntap1$1_0.well.n2 6.9865
R667 nmos_diode_2/ntap1$1_0.well.n2 nmos_diode_2/ntap1$1_0.well.t0 6.74476
R668 nmos_diode_2/ntap1$1_0.well.n3 nmos_diode_2/ntap1$1_0.well.t3 2.2081
R669 nmos_diode_2/ntap1$1_1.well nmos_diode_2/ntap1$1_0.well.n0 2.35302
R670 nmos_diode_2/ntap1$1_0.well.n3 nmos_diode_2/ntap1$1_0.well.n1 0.275228
R671 ena.n1 ena 32.2644
R672 ena.n4 ena.n3 10.0428
R673 ena.n3 ena.n2 9.01438
R674 ena.n1 ena.n0 9.00695
R675 ena.n0 ena.t2 7.51188
R676 ena.n2 ena.t1 7.50446
R677 ena.n4 ena.t0 2.11116
R678 ena.n3 ena.n1 0.8233
R679 ena ena.n4 0.292935
R680 ena.n2 ena 0.0470511
R681 ena.n0 ena 0.0396353
R682 ua[0].t1 ua[0].t0 40.8997
R683 ua[0] ua[0].t1 7.19763
R684 sg13g2_and2_2_1.X sg13g2_and2_2_1.X.t2 60.8893
R685 sg13g2_and2_2_1.X sg13g2_and2_2_1.X.t0 9.02833
R686 sg13g2_and2_2_1.X sg13g2_and2_2_1.X.t1 5.7736
C0 ua[0] uo_out[7] 49.64579f
C1 VPWR uo_out[7] 17.86373f
C2 sg13g2_and2_2_0.X uo_out[7] 18.47608f
C3 sg13g2_and2_2_1.X.t2 uo_out[7] 50.6667f
C4 nmos_diode_2/ntap1$1_0.well.t4 uo_out[7] 40.3662f
C5 nmos_diode_3/ntap1$1_0.well.t3 uo_out[7] 40.5949f
C6 nmos_diode_1/ntap1$1_0.well.t4 uo_out[7] 38.5116f
C7 sg13g2_and2_2_0.X.t2 uo_out[7] 43.8883f
C8 sg13g2_and2_2_0.X.t3 uo_out[7] 43.6818f
.ends

