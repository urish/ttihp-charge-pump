* Dickson Charge Pump Teshbench
* Run with `make sim`

.include "pdk_lib.spice"

.param temp=27
.param mc_ok = 1

* Power supply
V1 VGND 0 0
V2 VPWR VGND 1.2
* Clock
V3 clk VGND PULSE(0 1.2 0 0 0 250n 500n)
* Enable
V4 VPWR ena 0

* Output load
R1 ua[0] VGND 7Meg

.include "tt_um_urish_dickson_pump.spice"

x1 VGND VPWR clk ena rst_n
+ VGND VGND VGND VGND VGND VGND VGND VGND
+ VGND VGND VGND VGND VGND VGND VGND VGND
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ ua[0] ua[1] ua[2] ua[3]
+ tt_um_urish_dickson_pump

.tran 1n 100u

.control
run
plot "ua[0]" clk
.endc
.end

.end
